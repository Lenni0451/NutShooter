module main

const (
	game_name           = 'Nut Shooter'
	assets_font_regular = $embed_file('assets/OpenSans-Regular.ttf', .zlib)
	assets_font_bold    = $embed_file('assets/OpenSans-Bold.ttf', .zlib)
)
