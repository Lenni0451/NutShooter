module main

const game_name = 'Nut Shooter'
const assets_font_regular = $embed_file('assets/OpenSans-Regular.ttf', .zlib)
const assets_font_bold = $embed_file('assets/OpenSans-Bold.ttf', .zlib)
